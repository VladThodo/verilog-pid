// 64 bytes memory block

module memory(
    input clk_in,
    input reset,
    input write_enable,
    input [5:0] addr,
    input [7:0] data);

    always @(posedge clk_in) begin
       
    end

endmodule
